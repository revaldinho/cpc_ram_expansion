// 
// t35_romboard netlist
// 
// netlister.py format
// 
// (c) Revaldinho, 2018
// 
//  
module t35_romboard ();

  // wire declarations
  supply0 VSS;
  supply1 VDD_EXT;
  supply1 VDD_CPC;
  supply1 VDD;

  wire Sound;  
  wire A15,A14,A13,A12,A11,A10,A9,A8,A7,A6,A5,A4,A3,A2,A1,A0 ;
  wire D7,D6,D5,D4,D3,D2,D1,D0 ;
  wire MREQ_B;  
  wire M1_B;
  wire RFSH_B;
  wire IOREQ_B;
  wire RD_B;
  wire WR_B;
  wire HALT_B;
  wire INT_B ;
  wire NMI_B ;
  wire BUSRQ_B;  
  wire BUSACK_B;
  wire READY;
  wire BUSRESET_B;
  wire RESET_B;
  wire ROMEN_B;
  wire ROMDIS ;
  wire RAMRD_B;
  wire RAMDIS;
  wire CURSOR;
  wire LPEN;
  wire EXP_B;
  wire CLK;

  wire romdis_pre;
  wire dout0,dout1,dout2,dout3,dout4,dout5,dout6,dout7;
  
  // 3 pin header with link to use either CPC or external 5V power for the board
  hdr1x03      L1 (
                   .p1(VDD_CPC),
                   .p2(VDD),
                   .p3(VDD_EXT)
                   );

  // 3 pin Tabbed power connector for external 5V power
  powerheader3   CONN0 (
                        .vdd1(VDD_EXT),
                        .vdd2(VDD_EXT),
                        .gnd(VSS)
                        );

  // Radial electolytic, one per board on the main 5V supply
  cap22uf         CAP22UF(.minus(VSS),.plus(VDD));

  // Amstrad CPC Edge Connector
  //
  // V1.01 Corrected upper and lower rows

  idc_hdr_50w  CONN1 (
                      .p50(Sound),   .p49(VSS),
                      .p48(A15),     .p47(A14),
                      .p46(A13),     .p45(A12),
                      .p44(A11),     .p43(A10),
                      .p42(A9),      .p41(A8)
                      .p40(A7),      .p39(A6),
                      .p38(A5),      .p37(A4),
                      .p36(A3),      .p35(A2),
                      .p34(A1),      .p33(A0),
                      .p32(D7),      .p31(D6)
                      .p30(D5),      .p29(D4),
                      .p28(D3),      .p27(D2),
                      .p26(D1),      .p25(D0),
                      .p24(VDD_CPC), .p23(MREQ_B),
                      .p22(M1_B),    .p21(RFSH_B),
                      .p20(IOREQ_B), .p19(RD_B),
                      .p18(WR_B),    .p17(HALT_B),
                      .p16(INT_B),   .p15(NMI_B),
                      .p14(BUSRQ_B), .p13(BUSACK_B),
                      .p12(READY),   .p11(BUSRESET_B),
                      .p10(RESET_B), .p9 (ROMEN_B),
                      .p8 (ROMDIS),  .p7 (RAMRD_B),
                      .p6 (RAMDIS),  .p5 (CURSOR),
                      .p4 (LPEN),    .p3 (EXP_B),
                      .p2 (VSS),     .p1 (CLK),
                      ) ;



  teensy35_noxpins    U0 (
                  .gnd(VSS),       .vin(VDD),
                  .b16(A8),        .agnd(VSS),
                  .b17(A9),        .vdd_3v3_250ma(),
                  .d0(A0),         .c2(dout2),
                  .a12(),          .c1(dout1),
                  .a13(),          .d6(A6),
                  .d7(A7),         .d5(A5),
                  .d4(A4),         .b2(WR_B),
                  .d2(A2),         .b3(RAMRD_B),
                  .d3(A3),         .b1(IOREQ_B),
                  .c3(dout3),      .b0(MREQ_B),
                  .c4(dout4),      .c0(dout0),
                  .c6(dout6),      .d1(A1),
                  .c7(dout7),      .c5(dout5),
                  .vdd_3v3(),      .gnd2(VSS),
                  .e26(),          .dac1(),
                  .a5(),           .dac0(),
                  .a14(),          .a17(),
                  .a15(),          .c11(),
                  .a16(),          .c10(),
                  .b18(A10),       .c9(READY),
                  .b19(A11),       .c8(romvalid),
                  .b10(RD_B),      .e25(),
                  .b11(CLK),       .e24(),

	                          .vusb(),         
	                                                           
	          .nc(),          .aref(),         
	          .a26(),         .a10(),          
	          .a25(),         .a11(),          
	          .gnd1(VSS),     .e11(),          
	          .gnd4(VSS),     .e10(),          
	          .gnd5(VSS),     .d11(),          
	                          .d15(D3),        
	                                                   
	          .a28(),         .d12(D0),        
	          .a29(),         .d13(D1),        
	          .a26(),         .d14(D2),        
	          .b20(A12),      .b5(M1_B),       
	          .b22(A14),      .b4(ROMEN_B),    
	          .b23(A15),      .d9(),           
	          .b21(A13),      .d8(),           
	          .gnd(VSS),      .vdd_3v3_1(),
                  .vdd_3v3_2(),    
                  
                  .reset(),
                  .prog(),
                  .gnd(),
                  .vdd_3v3_2(),
                  .vbat()
                  );

  SN74245  U1 (
               .dir(VDD),     .vdd(VDD),
               .a0(D7),       .gb(bufoe_b),
               .a1(D6),       .b0(dout7),
               .a2(D5),       .b1(dout6),
               .a3(D4),       .b2(dout5),
               .a4(D3),       .b3(dout4),
               .a5(D2),       .b4(dout3),
               .a6(D1),       .b5(dout2),
               .a7(D0),       .b6(dout1),
               .vss(VSS),     .b7(dout0),
               );
  
  SN7400   U2 ( .i0_0(romvalid), .i0_1(A14), .o0(romdis_b),
                .i1_0(romdis_b), .i1_1(romdis_b), .o1(romdis_pre),
                .i2_0(ROMEN_B), .i2_1(ROMEN_B), .o2(romen),
                .i3_0(romen), .i3_1(romdis_pre), .o3(bufoe_b),
                .vss(VSS), .vdd(VDD)
               );
  
  
  DIODE_1N4148 D0 (
                .A(romdis_pre),
                .C(ROMDIS)
                );

   // Decoupling caps for 74 logic only - T35 has its own
   cap100nf CAP100N_1 (.p0( VSS ), .p1( VDD ));
   cap100nf CAP100N_2 (.p0( VSS ), .p1( VDD ));

endmodule
